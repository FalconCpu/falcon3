`timescale 1ns / 1ps

module sdram_arbiter(
    input clock,
    input reset,

    // Connections to the SDRAM controller
    output  logic [2:0]  sdram_req,          // Which bus master requests SDRAM access
    output  logic [25:0] sdram_addr,         // Address of data to read/write
    output  logic        sdram_write,        // 1 = write, 0 = read
    output  logic        sdram_burst,        // 1 = burst, 0 = single
    output  logic [3:0]  sdram_byte_enable,  // For a write, which bytes to write.
    output  logic [31:0] sdram_wdata,        // Data to write
    input   logic        sdram_ack,          // SDRAM has recieved the request (signal master to deassert)
    input   logic [31:0] sdram_rdata,        // Data read from SDRAM
    input   logic [2:0]  sdram_rdvalid,      // Which bus master the data is for
    input   logic        sdram_complete,     // SDRAM controller is done with the current burst

    // Bus master 1
    input   logic        bus1_request,
    input   logic [25:0] bus1_addr,
    input   logic        bus1_write,
    input   logic        bus1_burst,
    input   logic [3:0]  bus1_byte_enable,
    input   logic [31:0] bus1_wdata,
    output  logic        bus1_ack,
    output  logic [31:0] bus1_rdata,
    output  logic        bus1_rdvalid,
    output  logic        bus1_complete,

    // Bus master 2
    input   logic        bus2_request,
    input   logic [25:0] bus2_addr,
    input   logic        bus2_write,
    input   logic        bus2_burst,
    input   logic [3:0]  bus2_byte_enable,
    input   logic [31:0] bus2_wdata,
    output  logic        bus2_ack,
    output  logic [31:0] bus2_rdata,
    output  logic        bus2_rdvalid,
    output  logic        bus2_complete,

    // Bus master 3
    input   logic        bus3_request,
    input   logic [25:0] bus3_addr,
    input   logic        bus3_write,
    input   logic        bus3_burst,
    input   logic [3:0]  bus3_byte_enable,
    input   logic [31:0] bus3_wdata,
    output  logic        bus3_ack,
    output  logic [31:0] bus3_rdata,
    output  logic        bus3_rdvalid,
    output  logic        bus3_complete,

    // Bus master 4
    input   logic        bus4_request,
    input   logic [25:0] bus4_addr,
    input   logic        bus4_write,
    input   logic        bus4_burst,
    input   logic [3:0]  bus4_byte_enable,
    input   logic [31:0] bus4_wdata,
    output  logic        bus4_ack,
    output  logic [31:0] bus4_rdata,
    output  logic        bus4_rdvalid,
    output  logic        bus4_complete,

    // Bus master 5
    input   logic        bus5_request,
    input   logic [25:0] bus5_addr,
    input   logic        bus5_write,
    input   logic        bus5_burst,
    input   logic [3:0]  bus5_byte_enable,
    input   logic [31:0] bus5_wdata,
    output  logic        bus5_ack,
    output  logic [31:0] bus5_rdata,
    output  logic        bus5_rdvalid,
    output  logic        bus5_complete


);

logic [2:0]  next_req;
logic [25:0] next_addr;
logic        next_write;
logic        next_burst;
logic [3:0]  next_byte_enable;
logic [31:0] next_wdata;

// synthesis translate_off
integer fh;
initial fh = $fopen("rtl_mem.log");
// synthesis translate_on


always_comb begin
    next_req = sdram_req;
    next_addr = sdram_addr;
    next_write = sdram_write;
    next_burst = sdram_burst;
    next_byte_enable = sdram_byte_enable;
    next_wdata = sdram_wdata;
    bus1_ack = 1'b0;
    bus2_ack = 1'b0;
    bus3_ack = 1'b0;
    bus4_ack = 1'b0;
    bus5_ack = 1'b0;

    if (sdram_req==3'b000) begin
        if (bus1_request) begin
            next_req = 3'h1;
            next_addr = bus1_addr;
            next_write = bus1_write;
            next_burst = bus1_burst;
            next_byte_enable = bus1_byte_enable;
            next_wdata = bus1_wdata;
            bus1_ack = 1'b1;
        end else if (bus2_request) begin
            next_req = 3'h2;
            next_addr = bus2_addr;
            next_write = bus2_write;
            next_burst = bus2_burst;
            next_byte_enable = bus2_byte_enable;
            next_wdata = bus2_wdata;
            bus2_ack = 1'b1;

        end else if (bus3_request) begin
            next_req = 3'h3;
            next_addr = bus3_addr;
            next_write = bus3_write;
            next_burst = bus3_burst;
            next_byte_enable = bus3_byte_enable;
            next_wdata = bus3_wdata;
            bus3_ack = 1'b1;
        end else if (bus4_request) begin
            next_req = 3'h4;
            next_addr = bus4_addr;
            next_write = bus4_write;
            next_burst = bus4_burst;
            next_byte_enable = bus4_byte_enable;
            next_wdata = bus4_wdata;
            bus4_ack = 1'b1;
        end else if (bus5_request) begin
            next_req = 3'h5;
            next_addr = bus5_addr;
            next_write = bus5_write;
            next_burst = bus5_burst;
            next_byte_enable = bus5_byte_enable;
            next_wdata = bus5_wdata;
            bus5_ack = 1'b1;
        end
    end

    if (sdram_ack) begin
        next_req = 3'b000;
        next_addr = 26'bx;
        next_write = 1'b0;
        next_burst = 1'b0;
        next_byte_enable = 4'bx;
        next_wdata = 32'bx;
    end

    // Pass data from the SDRAM controller to the bus master
    bus1_rdata = (sdram_rdvalid==3'h1) ? sdram_rdata : 32'bx;
    bus2_rdata = (sdram_rdvalid==3'h2) ? sdram_rdata : 32'bx;
    bus3_rdata = (sdram_rdvalid==3'h3) ? sdram_rdata : 32'bx;
    bus4_rdata = (sdram_rdvalid==3'h4) ? sdram_rdata : 32'bx;
    bus5_rdata = (sdram_rdvalid==3'h5) ? sdram_rdata : 32'bx;
    bus1_rdvalid = sdram_rdvalid==3'h1;
    bus2_rdvalid = sdram_rdvalid==3'h2;
    bus3_rdvalid = sdram_rdvalid==3'h3;
    bus4_rdvalid = sdram_rdvalid==3'h4;
    bus5_rdvalid = sdram_rdvalid==3'h5;
    bus1_complete = sdram_complete && sdram_rdvalid==3'h1;
    bus2_complete = sdram_complete && sdram_rdvalid==3'h2;
    bus3_complete = sdram_complete && sdram_rdvalid==3'h3;
    bus4_complete = sdram_complete && sdram_rdvalid==3'h4;
    bus5_complete = sdram_complete && sdram_rdvalid==3'h5;

    if (reset) begin
        next_req = 3'b000;
    end
end

always_ff @(posedge clock) begin
    sdram_req <= next_req;
    sdram_addr <= next_addr;
    sdram_write <= next_write;
    sdram_burst <= next_burst;
    sdram_byte_enable <= next_byte_enable;
    sdram_wdata <= next_wdata;

    // synthesis translate_off
    if (sdram_req == 3'b000 && sdram_ack)
        $display("Error: %t SDRAM arbiter received ack without a request", $time);

    if (sdram_req==3'h0 && next_req==3'h2 && bus2_write)
        $fwrite(fh, "[%08x]=%08x %x\n", bus2_addr, bus2_wdata, bus2_byte_enable);
    // synthesis translate_on


end

endmodule